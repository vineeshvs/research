// Full Adder rtl

module full_adder (a0, b0, c0, a1, b1, c_out, s_out, s2, s3);

   // Inputs_top
   // Outputs_top

output d1
output c3